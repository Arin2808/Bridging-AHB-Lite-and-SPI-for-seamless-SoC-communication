package fifo_pkg;
    import uvm_pkg::*;
`include "fifo_transaction.sv"
`include "fifo_sequence.sv"
`include "fifo_driver.sv"
`include "fifo_monitor.sv"
`include "fifo_scoreboard.sv"
`include "fifo_agent.sv"
`include "fifo_env.sv"
`include "fifo_test.sv"
// `include "fifo_if.sv"
endpackage